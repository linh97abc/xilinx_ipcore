
`timescale 1 ns / 1 ps

	module axi_fifo_uart_v1_0 #
	(
		// Users to add parameters here
        parameter integer C_S00_AXI_CLK_FREQ_HZ = 100000000,
        parameter integer C_BAUDRATE     = 115200,
        parameter integer C_PARITY = 0, 			/* 0(none), 1(even), 2(odd), 3(mark), 4(space) */
        parameter integer C_DATA_BITS = 8, 		/* Byte Size (16 max) */
        parameter integer C_STOP_BITS = 0, 		/* 0(one stop), 1(two stops) */
        parameter integer C_FIFO_DEPTH = 256,		/* FIFO Depth */
		// User parameters ends
		// Do not modify the parameters beyond this line


		// Parameters of Axi Slave Bus Interface S00_AXI
		parameter integer C_S00_AXI_DATA_WIDTH	= 32,
		parameter integer C_S00_AXI_ADDR_WIDTH	= 6
	)
	(
		// Users to add ports here
		output irq,
	   // UART Port
        output wire tx,
        input wire rx,
        
		// User ports ends
		// Do not modify the ports beyond this line


		// Ports of Axi Slave Bus Interface S00_AXI
		input wire  s00_axi_aclk,
		input wire  s00_axi_aresetn,
		input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_awaddr,
		input wire [2 : 0] s00_axi_awprot,
		input wire  s00_axi_awvalid,
		output wire  s00_axi_awready,
		input wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_wdata,
		input wire [(C_S00_AXI_DATA_WIDTH/8)-1 : 0] s00_axi_wstrb,
		input wire  s00_axi_wvalid,
		output wire  s00_axi_wready,
		output wire [1 : 0] s00_axi_bresp,
		output wire  s00_axi_bvalid,
		input wire  s00_axi_bready,
		input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_araddr,
		input wire [2 : 0] s00_axi_arprot,
		input wire  s00_axi_arvalid,
		output wire  s00_axi_arready,
		output wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_rdata,
		output wire [1 : 0] s00_axi_rresp,
		output wire  s00_axi_rvalid,
		input wire  s00_axi_rready
	);
// Instantiation of Axi Bus Interface S00_AXI
	axi_fifo_uart_v1_0_S00_AXI # ( 
        .ACLK_FREQ_HZ(C_S00_AXI_CLK_FREQ_HZ),
        .BAUDRATE(C_BAUDRATE),
        .PARITY(C_PARITY), 			/* 0(none), 1(even), 2(odd), 3(mark), 4(space) */
        .BYTE_SIZE(C_DATA_BITS), 		/* Byte Size (16 max) */
        .STOP_BITS(C_STOP_BITS), 		/* 0(one stop), 1(two stops) */
        .FIFO_DEPTH(C_FIFO_DEPTH),		/* FIFO Depth */
        //
		.C_S_AXI_DATA_WIDTH(C_S00_AXI_DATA_WIDTH),
		.C_S_AXI_ADDR_WIDTH(C_S00_AXI_ADDR_WIDTH)
	) axi_fifo_uart_v1_0_S00_AXI_inst (
        .irq(irq),
        .tx(tx),
        .rx(rx),
        //
		.S_AXI_ACLK(s00_axi_aclk),
		.S_AXI_ARESETN(s00_axi_aresetn),
		.S_AXI_AWADDR(s00_axi_awaddr),
		.S_AXI_AWPROT(s00_axi_awprot),
		.S_AXI_AWVALID(s00_axi_awvalid),
		.S_AXI_AWREADY(s00_axi_awready),
		.S_AXI_WDATA(s00_axi_wdata),
		.S_AXI_WSTRB(s00_axi_wstrb),
		.S_AXI_WVALID(s00_axi_wvalid),
		.S_AXI_WREADY(s00_axi_wready),
		.S_AXI_BRESP(s00_axi_bresp),
		.S_AXI_BVALID(s00_axi_bvalid),
		.S_AXI_BREADY(s00_axi_bready),
		.S_AXI_ARADDR(s00_axi_araddr),
		.S_AXI_ARPROT(s00_axi_arprot),
		.S_AXI_ARVALID(s00_axi_arvalid),
		.S_AXI_ARREADY(s00_axi_arready),
		.S_AXI_RDATA(s00_axi_rdata),
		.S_AXI_RRESP(s00_axi_rresp),
		.S_AXI_RVALID(s00_axi_rvalid),
		.S_AXI_RREADY(s00_axi_rready)
	);

	// Add user logic here

	// User logic ends

	endmodule
